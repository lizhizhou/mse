// qsys.v

// Generated using ACDS version 12.1sp1 243 at 2013.08.05.09:56:08

`timescale 1 ps / 1 ps
module qsys (
		inout  wire  port1_P0,               //            port1.P0
		inout  wire  port1_P1,               //                 .P1
		inout  wire  port1_P2,               //                 .P2
		inout  wire  port1_P3,               //                 .P3
		inout  wire  port1_P4,               //                 .P4
		inout  wire  port1_P5,               //                 .P5
		inout  wire  port1_P6,               //                 .P6
		inout  wire  port1_P7,               //                 .P7
		output wire  led_export,             //              led.export
		output wire  dryer_export,           //            dryer.export
		output wire  qsys_serial_host_sdo,   // qsys_serial_host.sdo
		input  wire  qsys_serial_host_sdi,   //                 .sdi
		input  wire  qsys_serial_host_clk,   //                 .clk
		input  wire  qsys_serial_host_sle,   //                 .sle
		output wire  qsys_serial_host_srdy,  //                 .srdy
		input  wire  qsys_serial_host_reset, //                 .reset
		output wire  humidifier_export,      //       humidifier.export
		output wire  semi_cooler_HX,         //      semi_cooler.HX
		output wire  semi_cooler_HY,         //                 .HY
		inout  wire  port0_P0,               //            port0.P0
		inout  wire  port0_P1,               //                 .P1
		inout  wire  port0_P2,               //                 .P2
		inout  wire  port0_P3,               //                 .P3
		inout  wire  port0_P4,               //                 .P4
		inout  wire  port0_P5,               //                 .P5
		inout  wire  port0_P6,               //                 .P6
		inout  wire  port0_P7,               //                 .P7
		output wire  humidifier_fan_export   //   humidifier_fan.export
	);

	wire         qsys_serial_host_0_mrst_reset;                                                                  // qsys_serial_host_0:rso_MRST_reset -> [PIO8_0:rsi_MRST_reset, PIO8_0_gpio_translator:reset, PIO8_0_gpio_translator_avalon_universal_slave_0_agent:reset, PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, PIO8_1:rsi_MRST_reset, PIO8_1_gpio_translator:reset, PIO8_1_gpio_translator_avalon_universal_slave_0_agent:reset, PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, brush_motor_driver_0:rsi_MRST_reset, brush_motor_driver_0:rsi_PWMRST_reset, brush_motor_driver_0_ctrl_translator:reset, brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:reset, brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, fan_motor_driver_0:rsi_MRST_reset, fan_motor_driver_0:rsi_PWMRST_reset, fan_motor_driver_0_ctrl_translator:reset, fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:reset, fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fan_motor_driver_1:rsi_MRST_reset, fan_motor_driver_1:rsi_PWMRST_reset, fan_motor_driver_1_ctrl_translator:reset, fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:reset, fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fan_motor_driver_2:rsi_MRST_reset, fan_motor_driver_2:rsi_PWMRST_reset, fan_motor_driver_2_ctrl_translator:reset, fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:reset, fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fan_motor_driver_3:rsi_MRST_reset, fan_motor_driver_3:rsi_PWMRST_reset, fan_motor_driver_3_ctrl_translator:reset, fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:reset, fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, limiter:reset, qsys_serial_host_0_m1_translator:reset, qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_mux:reset]
	wire         qsys_serial_host_0_mclk_clk;                                                                    // qsys_serial_host_0:cso_MCLK_clk -> [PIO8_0:csi_MCLK_clk, PIO8_0_gpio_translator:clk, PIO8_0_gpio_translator_avalon_universal_slave_0_agent:clk, PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, PIO8_1:csi_MCLK_clk, PIO8_1_gpio_translator:clk, PIO8_1_gpio_translator_avalon_universal_slave_0_agent:clk, PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, brush_motor_driver_0:csi_MCLK_clk, brush_motor_driver_0:csi_PWMCLK_clk, brush_motor_driver_0_ctrl_translator:clk, brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:clk, brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, fan_motor_driver_0:csi_MCLK_clk, fan_motor_driver_0:csi_PWMCLK_clk, fan_motor_driver_0_ctrl_translator:clk, fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:clk, fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, fan_motor_driver_1:csi_MCLK_clk, fan_motor_driver_1:csi_PWMCLK_clk, fan_motor_driver_1_ctrl_translator:clk, fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:clk, fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, fan_motor_driver_2:csi_MCLK_clk, fan_motor_driver_2:csi_PWMCLK_clk, fan_motor_driver_2_ctrl_translator:clk, fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:clk, fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, fan_motor_driver_3:csi_MCLK_clk, fan_motor_driver_3:csi_PWMCLK_clk, fan_motor_driver_3_ctrl_translator:clk, fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:clk, fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, limiter:clk, qsys_serial_host_0_m1_translator:clk, qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_mux:clk]
	wire         qsys_serial_host_0_m1_waitrequest;                                                              // qsys_serial_host_0_m1_translator:av_waitrequest -> qsys_serial_host_0:avm_M1_waitrequest
	wire   [7:0] qsys_serial_host_0_m1_address;                                                                  // qsys_serial_host_0:avm_M1_address -> qsys_serial_host_0_m1_translator:av_address
	wire  [31:0] qsys_serial_host_0_m1_writedata;                                                                // qsys_serial_host_0:avm_M1_writedata -> qsys_serial_host_0_m1_translator:av_writedata
	wire         qsys_serial_host_0_m1_write;                                                                    // qsys_serial_host_0:avm_M1_write -> qsys_serial_host_0_m1_translator:av_write
	wire         qsys_serial_host_0_m1_read;                                                                     // qsys_serial_host_0:avm_M1_read -> qsys_serial_host_0_m1_translator:av_read
	wire  [31:0] qsys_serial_host_0_m1_readdata;                                                                 // qsys_serial_host_0_m1_translator:av_readdata -> qsys_serial_host_0:avm_M1_readdata
	wire         qsys_serial_host_0_m1_begintransfer;                                                            // qsys_serial_host_0:avm_M1_begintransfer -> qsys_serial_host_0_m1_translator:av_begintransfer
	wire         qsys_serial_host_0_m1_readdatavalid;                                                            // qsys_serial_host_0_m1_translator:av_readdatavalid -> qsys_serial_host_0:avm_M1_readdatavalid
	wire   [3:0] qsys_serial_host_0_m1_byteenable;                                                               // qsys_serial_host_0:avm_M1_byteenable -> qsys_serial_host_0_m1_translator:av_byteenable
	wire         pio8_0_gpio_translator_avalon_anti_slave_0_waitrequest;                                         // PIO8_0:avs_gpio_waitrequest -> PIO8_0_gpio_translator:av_waitrequest
	wire  [31:0] pio8_0_gpio_translator_avalon_anti_slave_0_writedata;                                           // PIO8_0_gpio_translator:av_writedata -> PIO8_0:avs_gpio_writedata
	wire   [2:0] pio8_0_gpio_translator_avalon_anti_slave_0_address;                                             // PIO8_0_gpio_translator:av_address -> PIO8_0:avs_gpio_address
	wire         pio8_0_gpio_translator_avalon_anti_slave_0_write;                                               // PIO8_0_gpio_translator:av_write -> PIO8_0:avs_gpio_write
	wire         pio8_0_gpio_translator_avalon_anti_slave_0_read;                                                // PIO8_0_gpio_translator:av_read -> PIO8_0:avs_gpio_read
	wire  [31:0] pio8_0_gpio_translator_avalon_anti_slave_0_readdata;                                            // PIO8_0:avs_gpio_readdata -> PIO8_0_gpio_translator:av_readdata
	wire   [3:0] pio8_0_gpio_translator_avalon_anti_slave_0_byteenable;                                          // PIO8_0_gpio_translator:av_byteenable -> PIO8_0:avs_gpio_byteenable
	wire         pio8_1_gpio_translator_avalon_anti_slave_0_waitrequest;                                         // PIO8_1:avs_gpio_waitrequest -> PIO8_1_gpio_translator:av_waitrequest
	wire  [31:0] pio8_1_gpio_translator_avalon_anti_slave_0_writedata;                                           // PIO8_1_gpio_translator:av_writedata -> PIO8_1:avs_gpio_writedata
	wire   [2:0] pio8_1_gpio_translator_avalon_anti_slave_0_address;                                             // PIO8_1_gpio_translator:av_address -> PIO8_1:avs_gpio_address
	wire         pio8_1_gpio_translator_avalon_anti_slave_0_write;                                               // PIO8_1_gpio_translator:av_write -> PIO8_1:avs_gpio_write
	wire         pio8_1_gpio_translator_avalon_anti_slave_0_read;                                                // PIO8_1_gpio_translator:av_read -> PIO8_1:avs_gpio_read
	wire  [31:0] pio8_1_gpio_translator_avalon_anti_slave_0_readdata;                                            // PIO8_1:avs_gpio_readdata -> PIO8_1_gpio_translator:av_readdata
	wire   [3:0] pio8_1_gpio_translator_avalon_anti_slave_0_byteenable;                                          // PIO8_1_gpio_translator:av_byteenable -> PIO8_1:avs_gpio_byteenable
	wire         fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_waitrequest;                             // fan_motor_driver_0:avs_ctrl_waitrequest -> fan_motor_driver_0_ctrl_translator:av_waitrequest
	wire  [31:0] fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_writedata;                               // fan_motor_driver_0_ctrl_translator:av_writedata -> fan_motor_driver_0:avs_ctrl_writedata
	wire   [2:0] fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_address;                                 // fan_motor_driver_0_ctrl_translator:av_address -> fan_motor_driver_0:avs_ctrl_address
	wire         fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_write;                                   // fan_motor_driver_0_ctrl_translator:av_write -> fan_motor_driver_0:avs_ctrl_write
	wire         fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_read;                                    // fan_motor_driver_0_ctrl_translator:av_read -> fan_motor_driver_0:avs_ctrl_read
	wire  [31:0] fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_readdata;                                // fan_motor_driver_0:avs_ctrl_readdata -> fan_motor_driver_0_ctrl_translator:av_readdata
	wire   [3:0] fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_byteenable;                              // fan_motor_driver_0_ctrl_translator:av_byteenable -> fan_motor_driver_0:avs_ctrl_byteenable
	wire         fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_waitrequest;                             // fan_motor_driver_1:avs_ctrl_waitrequest -> fan_motor_driver_1_ctrl_translator:av_waitrequest
	wire  [31:0] fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_writedata;                               // fan_motor_driver_1_ctrl_translator:av_writedata -> fan_motor_driver_1:avs_ctrl_writedata
	wire   [2:0] fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_address;                                 // fan_motor_driver_1_ctrl_translator:av_address -> fan_motor_driver_1:avs_ctrl_address
	wire         fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_write;                                   // fan_motor_driver_1_ctrl_translator:av_write -> fan_motor_driver_1:avs_ctrl_write
	wire         fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_read;                                    // fan_motor_driver_1_ctrl_translator:av_read -> fan_motor_driver_1:avs_ctrl_read
	wire  [31:0] fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_readdata;                                // fan_motor_driver_1:avs_ctrl_readdata -> fan_motor_driver_1_ctrl_translator:av_readdata
	wire   [3:0] fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_byteenable;                              // fan_motor_driver_1_ctrl_translator:av_byteenable -> fan_motor_driver_1:avs_ctrl_byteenable
	wire         fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_waitrequest;                             // fan_motor_driver_2:avs_ctrl_waitrequest -> fan_motor_driver_2_ctrl_translator:av_waitrequest
	wire  [31:0] fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_writedata;                               // fan_motor_driver_2_ctrl_translator:av_writedata -> fan_motor_driver_2:avs_ctrl_writedata
	wire   [2:0] fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_address;                                 // fan_motor_driver_2_ctrl_translator:av_address -> fan_motor_driver_2:avs_ctrl_address
	wire         fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_write;                                   // fan_motor_driver_2_ctrl_translator:av_write -> fan_motor_driver_2:avs_ctrl_write
	wire         fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_read;                                    // fan_motor_driver_2_ctrl_translator:av_read -> fan_motor_driver_2:avs_ctrl_read
	wire  [31:0] fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_readdata;                                // fan_motor_driver_2:avs_ctrl_readdata -> fan_motor_driver_2_ctrl_translator:av_readdata
	wire   [3:0] fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_byteenable;                              // fan_motor_driver_2_ctrl_translator:av_byteenable -> fan_motor_driver_2:avs_ctrl_byteenable
	wire         brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // brush_motor_driver_0:avs_ctrl_waitrequest -> brush_motor_driver_0_ctrl_translator:av_waitrequest
	wire  [31:0] brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_writedata;                             // brush_motor_driver_0_ctrl_translator:av_writedata -> brush_motor_driver_0:avs_ctrl_writedata
	wire   [2:0] brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_address;                               // brush_motor_driver_0_ctrl_translator:av_address -> brush_motor_driver_0:avs_ctrl_address
	wire         brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_write;                                 // brush_motor_driver_0_ctrl_translator:av_write -> brush_motor_driver_0:avs_ctrl_write
	wire         brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_read;                                  // brush_motor_driver_0_ctrl_translator:av_read -> brush_motor_driver_0:avs_ctrl_read
	wire  [31:0] brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_readdata;                              // brush_motor_driver_0:avs_ctrl_readdata -> brush_motor_driver_0_ctrl_translator:av_readdata
	wire   [3:0] brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_byteenable;                            // brush_motor_driver_0_ctrl_translator:av_byteenable -> brush_motor_driver_0:avs_ctrl_byteenable
	wire         fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_waitrequest;                             // fan_motor_driver_3:avs_ctrl_waitrequest -> fan_motor_driver_3_ctrl_translator:av_waitrequest
	wire  [31:0] fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_writedata;                               // fan_motor_driver_3_ctrl_translator:av_writedata -> fan_motor_driver_3:avs_ctrl_writedata
	wire   [2:0] fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_address;                                 // fan_motor_driver_3_ctrl_translator:av_address -> fan_motor_driver_3:avs_ctrl_address
	wire         fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_write;                                   // fan_motor_driver_3_ctrl_translator:av_write -> fan_motor_driver_3:avs_ctrl_write
	wire         fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_read;                                    // fan_motor_driver_3_ctrl_translator:av_read -> fan_motor_driver_3:avs_ctrl_read
	wire  [31:0] fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_readdata;                                // fan_motor_driver_3:avs_ctrl_readdata -> fan_motor_driver_3_ctrl_translator:av_readdata
	wire   [3:0] fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_byteenable;                              // fan_motor_driver_3_ctrl_translator:av_byteenable -> fan_motor_driver_3:avs_ctrl_byteenable
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest;                         // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_waitrequest -> qsys_serial_host_0_m1_translator:uav_waitrequest
	wire   [2:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount;                          // qsys_serial_host_0_m1_translator:uav_burstcount -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata;                           // qsys_serial_host_0_m1_translator:uav_writedata -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_writedata
	wire   [9:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_address;                             // qsys_serial_host_0_m1_translator:uav_address -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_address
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock;                                // qsys_serial_host_0_m1_translator:uav_lock -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_lock
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_write;                               // qsys_serial_host_0_m1_translator:uav_write -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_write
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_read;                                // qsys_serial_host_0_m1_translator:uav_read -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata;                            // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_readdata -> qsys_serial_host_0_m1_translator:uav_readdata
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess;                         // qsys_serial_host_0_m1_translator:uav_debugaccess -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable;                          // qsys_serial_host_0_m1_translator:uav_byteenable -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_byteenable
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid;                       // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:av_readdatavalid -> qsys_serial_host_0_m1_translator:uav_readdatavalid
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // PIO8_0_gpio_translator:uav_waitrequest -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_burstcount -> PIO8_0_gpio_translator:uav_burstcount
	wire  [31:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_writedata;                             // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_writedata -> PIO8_0_gpio_translator:uav_writedata
	wire   [9:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_address;                               // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_address -> PIO8_0_gpio_translator:uav_address
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_write;                                 // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_write -> PIO8_0_gpio_translator:uav_write
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_lock;                                  // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_lock -> PIO8_0_gpio_translator:uav_lock
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_read;                                  // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_read -> PIO8_0_gpio_translator:uav_read
	wire  [31:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_readdata;                              // PIO8_0_gpio_translator:uav_readdata -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // PIO8_0_gpio_translator:uav_readdatavalid -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PIO8_0_gpio_translator:uav_debugaccess
	wire   [3:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:m0_byteenable -> PIO8_0_gpio_translator:uav_byteenable
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_source_valid -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_data;                           // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_source_data -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // PIO8_1_gpio_translator:uav_waitrequest -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_burstcount -> PIO8_1_gpio_translator:uav_burstcount
	wire  [31:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_writedata;                             // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_writedata -> PIO8_1_gpio_translator:uav_writedata
	wire   [9:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_address;                               // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_address -> PIO8_1_gpio_translator:uav_address
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_write;                                 // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_write -> PIO8_1_gpio_translator:uav_write
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_lock;                                  // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_lock -> PIO8_1_gpio_translator:uav_lock
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_read;                                  // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_read -> PIO8_1_gpio_translator:uav_read
	wire  [31:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_readdata;                              // PIO8_1_gpio_translator:uav_readdata -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // PIO8_1_gpio_translator:uav_readdatavalid -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_debugaccess -> PIO8_1_gpio_translator:uav_debugaccess
	wire   [3:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:m0_byteenable -> PIO8_1_gpio_translator:uav_byteenable
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_source_valid -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_data;                           // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_source_data -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rf_sink_ready -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // fan_motor_driver_0_ctrl_translator:uav_waitrequest -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;                // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> fan_motor_driver_0_ctrl_translator:uav_burstcount
	wire  [31:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                 // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> fan_motor_driver_0_ctrl_translator:uav_writedata
	wire   [9:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                   // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> fan_motor_driver_0_ctrl_translator:uav_address
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                     // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> fan_motor_driver_0_ctrl_translator:uav_write
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                      // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> fan_motor_driver_0_ctrl_translator:uav_lock
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                      // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> fan_motor_driver_0_ctrl_translator:uav_read
	wire  [31:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                  // fan_motor_driver_0_ctrl_translator:uav_readdata -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // fan_motor_driver_0_ctrl_translator:uav_readdatavalid -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fan_motor_driver_0_ctrl_translator:uav_debugaccess
	wire   [3:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;                // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> fan_motor_driver_0_ctrl_translator:uav_byteenable
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;              // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;               // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;              // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // fan_motor_driver_1_ctrl_translator:uav_waitrequest -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;                // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> fan_motor_driver_1_ctrl_translator:uav_burstcount
	wire  [31:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                 // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> fan_motor_driver_1_ctrl_translator:uav_writedata
	wire   [9:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                   // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> fan_motor_driver_1_ctrl_translator:uav_address
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                     // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> fan_motor_driver_1_ctrl_translator:uav_write
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                      // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> fan_motor_driver_1_ctrl_translator:uav_lock
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                      // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> fan_motor_driver_1_ctrl_translator:uav_read
	wire  [31:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                  // fan_motor_driver_1_ctrl_translator:uav_readdata -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // fan_motor_driver_1_ctrl_translator:uav_readdatavalid -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fan_motor_driver_1_ctrl_translator:uav_debugaccess
	wire   [3:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;                // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> fan_motor_driver_1_ctrl_translator:uav_byteenable
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;              // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;               // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;              // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // fan_motor_driver_2_ctrl_translator:uav_waitrequest -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;                // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> fan_motor_driver_2_ctrl_translator:uav_burstcount
	wire  [31:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                 // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> fan_motor_driver_2_ctrl_translator:uav_writedata
	wire   [9:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                   // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> fan_motor_driver_2_ctrl_translator:uav_address
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                     // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> fan_motor_driver_2_ctrl_translator:uav_write
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                      // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> fan_motor_driver_2_ctrl_translator:uav_lock
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                      // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> fan_motor_driver_2_ctrl_translator:uav_read
	wire  [31:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                  // fan_motor_driver_2_ctrl_translator:uav_readdata -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // fan_motor_driver_2_ctrl_translator:uav_readdatavalid -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fan_motor_driver_2_ctrl_translator:uav_debugaccess
	wire   [3:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;                // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> fan_motor_driver_2_ctrl_translator:uav_byteenable
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;              // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;               // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;              // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // brush_motor_driver_0_ctrl_translator:uav_waitrequest -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> brush_motor_driver_0_ctrl_translator:uav_burstcount
	wire  [31:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> brush_motor_driver_0_ctrl_translator:uav_writedata
	wire   [9:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> brush_motor_driver_0_ctrl_translator:uav_address
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> brush_motor_driver_0_ctrl_translator:uav_write
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> brush_motor_driver_0_ctrl_translator:uav_lock
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> brush_motor_driver_0_ctrl_translator:uav_read
	wire  [31:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // brush_motor_driver_0_ctrl_translator:uav_readdata -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // brush_motor_driver_0_ctrl_translator:uav_readdatavalid -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> brush_motor_driver_0_ctrl_translator:uav_debugaccess
	wire   [3:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> brush_motor_driver_0_ctrl_translator:uav_byteenable
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // fan_motor_driver_3_ctrl_translator:uav_waitrequest -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;                // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> fan_motor_driver_3_ctrl_translator:uav_burstcount
	wire  [31:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                 // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> fan_motor_driver_3_ctrl_translator:uav_writedata
	wire   [9:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                   // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> fan_motor_driver_3_ctrl_translator:uav_address
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                     // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> fan_motor_driver_3_ctrl_translator:uav_write
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                      // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> fan_motor_driver_3_ctrl_translator:uav_lock
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                      // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> fan_motor_driver_3_ctrl_translator:uav_read
	wire  [31:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                  // fan_motor_driver_3_ctrl_translator:uav_readdata -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // fan_motor_driver_3_ctrl_translator:uav_readdatavalid -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fan_motor_driver_3_ctrl_translator:uav_debugaccess
	wire   [3:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;                // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> fan_motor_driver_3_ctrl_translator:uav_byteenable
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;              // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;               // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;              // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_endofpacket;                // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_valid;                      // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_startofpacket;              // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [82:0] qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_data;                       // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router:sink_ready -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:cp_ready
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_valid;                                 // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [82:0] pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_data;                                  // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router:sink_ready -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_valid;                                 // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [82:0] pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_data;                                  // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_001:sink_ready -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                     // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [82:0] fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                      // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_002:sink_ready -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                     // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [82:0] fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                      // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_003:sink_ready -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                     // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [82:0] fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                      // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_004:sink_ready -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [82:0] brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                     // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [82:0] fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                      // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_006:sink_ready -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                    // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                          // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                  // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [82:0] addr_router_src_data;                                                                           // addr_router:src_data -> limiter:cmd_sink_data
	wire   [6:0] addr_router_src_channel;                                                                        // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                          // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                    // limiter:rsp_src_endofpacket -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                          // limiter:rsp_src_valid -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                  // limiter:rsp_src_startofpacket -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [82:0] limiter_rsp_src_data;                                                                           // limiter:rsp_src_data -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_data
	wire   [6:0] limiter_rsp_src_channel;                                                                        // limiter:rsp_src_channel -> qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                          // qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                                // cmd_xbar_demux:src0_endofpacket -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                      // cmd_xbar_demux:src0_valid -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                              // cmd_xbar_demux:src0_startofpacket -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src0_data;                                                                       // cmd_xbar_demux:src0_data -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src0_channel;                                                                    // cmd_xbar_demux:src0_channel -> PIO8_0_gpio_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src1_endofpacket;                                                                // cmd_xbar_demux:src1_endofpacket -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                      // cmd_xbar_demux:src1_valid -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                              // cmd_xbar_demux:src1_startofpacket -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src1_data;                                                                       // cmd_xbar_demux:src1_data -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src1_channel;                                                                    // cmd_xbar_demux:src1_channel -> PIO8_1_gpio_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src2_endofpacket;                                                                // cmd_xbar_demux:src2_endofpacket -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                      // cmd_xbar_demux:src2_valid -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                              // cmd_xbar_demux:src2_startofpacket -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src2_data;                                                                       // cmd_xbar_demux:src2_data -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src2_channel;                                                                    // cmd_xbar_demux:src2_channel -> fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src3_endofpacket;                                                                // cmd_xbar_demux:src3_endofpacket -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                      // cmd_xbar_demux:src3_valid -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                              // cmd_xbar_demux:src3_startofpacket -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src3_data;                                                                       // cmd_xbar_demux:src3_data -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src3_channel;                                                                    // cmd_xbar_demux:src3_channel -> fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src4_endofpacket;                                                                // cmd_xbar_demux:src4_endofpacket -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                      // cmd_xbar_demux:src4_valid -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                              // cmd_xbar_demux:src4_startofpacket -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src4_data;                                                                       // cmd_xbar_demux:src4_data -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src4_channel;                                                                    // cmd_xbar_demux:src4_channel -> fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src5_endofpacket;                                                                // cmd_xbar_demux:src5_endofpacket -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                                      // cmd_xbar_demux:src5_valid -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                              // cmd_xbar_demux:src5_startofpacket -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src5_data;                                                                       // cmd_xbar_demux:src5_data -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src5_channel;                                                                    // cmd_xbar_demux:src5_channel -> brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src6_endofpacket;                                                                // cmd_xbar_demux:src6_endofpacket -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                                      // cmd_xbar_demux:src6_valid -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                              // cmd_xbar_demux:src6_startofpacket -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src6_data;                                                                       // cmd_xbar_demux:src6_data -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src6_channel;                                                                    // cmd_xbar_demux:src6_channel -> fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                      // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                              // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [82:0] rsp_xbar_demux_src0_data;                                                                       // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [6:0] rsp_xbar_demux_src0_channel;                                                                    // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                      // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                            // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                  // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                          // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [82:0] rsp_xbar_demux_001_src0_data;                                                                   // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [6:0] rsp_xbar_demux_001_src0_channel;                                                                // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                  // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                            // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                  // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                          // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [82:0] rsp_xbar_demux_002_src0_data;                                                                   // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [6:0] rsp_xbar_demux_002_src0_channel;                                                                // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                  // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                            // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                  // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                          // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [82:0] rsp_xbar_demux_003_src0_data;                                                                   // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [6:0] rsp_xbar_demux_003_src0_channel;                                                                // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                  // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                            // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                  // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                          // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [82:0] rsp_xbar_demux_004_src0_data;                                                                   // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [6:0] rsp_xbar_demux_004_src0_channel;                                                                // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                  // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                            // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                  // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                          // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [82:0] rsp_xbar_demux_005_src0_data;                                                                   // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [6:0] rsp_xbar_demux_005_src0_channel;                                                                // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                  // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                            // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                  // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                          // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [82:0] rsp_xbar_demux_006_src0_data;                                                                   // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [6:0] rsp_xbar_demux_006_src0_channel;                                                                // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                  // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                    // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                  // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [82:0] limiter_cmd_src_data;                                                                           // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [6:0] limiter_cmd_src_channel;                                                                        // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                          // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                   // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                         // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                 // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [82:0] rsp_xbar_mux_src_data;                                                                          // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [6:0] rsp_xbar_mux_src_channel;                                                                       // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                         // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         cmd_xbar_demux_src0_ready;                                                                      // PIO8_0_gpio_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                                      // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                            // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                    // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [82:0] id_router_src_data;                                                                             // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [6:0] id_router_src_channel;                                                                          // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                            // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                                      // PIO8_1_gpio_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                                  // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                        // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [82:0] id_router_001_src_data;                                                                         // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [6:0] id_router_001_src_channel;                                                                      // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                        // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_src2_ready;                                                                      // fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire         id_router_002_src_endofpacket;                                                                  // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                        // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [82:0] id_router_002_src_data;                                                                         // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [6:0] id_router_002_src_channel;                                                                      // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                        // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_src3_ready;                                                                      // fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire         id_router_003_src_endofpacket;                                                                  // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                        // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [82:0] id_router_003_src_data;                                                                         // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [6:0] id_router_003_src_channel;                                                                      // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                        // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_src4_ready;                                                                      // fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src4_ready
	wire         id_router_004_src_endofpacket;                                                                  // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                        // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [82:0] id_router_004_src_data;                                                                         // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [6:0] id_router_004_src_channel;                                                                      // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                        // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_src5_ready;                                                                      // brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src5_ready
	wire         id_router_005_src_endofpacket;                                                                  // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                        // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [82:0] id_router_005_src_data;                                                                         // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [6:0] id_router_005_src_channel;                                                                      // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                        // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_src6_ready;                                                                      // fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src6_ready
	wire         id_router_006_src_endofpacket;                                                                  // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                        // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [82:0] id_router_006_src_data;                                                                         // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [6:0] id_router_006_src_channel;                                                                      // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                        // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire   [6:0] limiter_cmd_valid_data;                                                                         // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid

	qsys_serial_host #(
		.initial_state (9'b000000000)
	) qsys_serial_host_0 (
		.rso_MRST_reset       (qsys_serial_host_0_mrst_reset),       //        mrst.reset
		.cso_MCLK_clk         (qsys_serial_host_0_mclk_clk),         //        mclk.clk
		.avm_M1_writedata     (qsys_serial_host_0_m1_writedata),     //          m1.writedata
		.avm_M1_readdata      (qsys_serial_host_0_m1_readdata),      //            .readdata
		.avm_M1_address       (qsys_serial_host_0_m1_address),       //            .address
		.avm_M1_byteenable    (qsys_serial_host_0_m1_byteenable),    //            .byteenable
		.avm_M1_write         (qsys_serial_host_0_m1_write),         //            .write
		.avm_M1_read          (qsys_serial_host_0_m1_read),          //            .read
		.avm_M1_begintransfer (qsys_serial_host_0_m1_begintransfer), //            .begintransfer
		.avm_M1_readdatavalid (qsys_serial_host_0_m1_readdatavalid), //            .readdatavalid
		.avm_M1_waitrequest   (qsys_serial_host_0_m1_waitrequest),   //            .waitrequest
		.sdo                  (qsys_serial_host_sdo),                // conduit_end.export
		.sdi                  (qsys_serial_host_sdi),                //            .export
		.clk                  (qsys_serial_host_clk),                //            .export
		.sle                  (qsys_serial_host_sle),                //            .export
		.srdy                 (qsys_serial_host_srdy),               //            .export
		.reset                (qsys_serial_host_reset)               //            .export
	);

	PIO8 pio8_0 (
		.rsi_MRST_reset       (qsys_serial_host_0_mrst_reset),                          // mrst.reset
		.csi_MCLK_clk         (qsys_serial_host_0_mclk_clk),                            // mclk.clk
		.avs_gpio_writedata   (pio8_0_gpio_translator_avalon_anti_slave_0_writedata),   // gpio.writedata
		.avs_gpio_readdata    (pio8_0_gpio_translator_avalon_anti_slave_0_readdata),    //     .readdata
		.avs_gpio_address     (pio8_0_gpio_translator_avalon_anti_slave_0_address),     //     .address
		.avs_gpio_byteenable  (pio8_0_gpio_translator_avalon_anti_slave_0_byteenable),  //     .byteenable
		.avs_gpio_write       (pio8_0_gpio_translator_avalon_anti_slave_0_write),       //     .write
		.avs_gpio_read        (pio8_0_gpio_translator_avalon_anti_slave_0_read),        //     .read
		.avs_gpio_waitrequest (pio8_0_gpio_translator_avalon_anti_slave_0_waitrequest), //     .waitrequest
		.coe_P0               (port0_P0),                                               //  PIO.export
		.coe_P1               (port0_P1),                                               //     .export
		.coe_P2               (port0_P2),                                               //     .export
		.coe_P3               (port0_P3),                                               //     .export
		.coe_P4               (port0_P4),                                               //     .export
		.coe_P5               (port0_P5),                                               //     .export
		.coe_P6               (port0_P6),                                               //     .export
		.coe_P7               (port0_P7)                                                //     .export
	);

	PIO8 pio8_1 (
		.rsi_MRST_reset       (qsys_serial_host_0_mrst_reset),                          // mrst.reset
		.csi_MCLK_clk         (qsys_serial_host_0_mclk_clk),                            // mclk.clk
		.avs_gpio_writedata   (pio8_1_gpio_translator_avalon_anti_slave_0_writedata),   // gpio.writedata
		.avs_gpio_readdata    (pio8_1_gpio_translator_avalon_anti_slave_0_readdata),    //     .readdata
		.avs_gpio_address     (pio8_1_gpio_translator_avalon_anti_slave_0_address),     //     .address
		.avs_gpio_byteenable  (pio8_1_gpio_translator_avalon_anti_slave_0_byteenable),  //     .byteenable
		.avs_gpio_write       (pio8_1_gpio_translator_avalon_anti_slave_0_write),       //     .write
		.avs_gpio_read        (pio8_1_gpio_translator_avalon_anti_slave_0_read),        //     .read
		.avs_gpio_waitrequest (pio8_1_gpio_translator_avalon_anti_slave_0_waitrequest), //     .waitrequest
		.coe_P0               (port1_P0),                                               //  PIO.export
		.coe_P1               (port1_P1),                                               //     .export
		.coe_P2               (port1_P2),                                               //     .export
		.coe_P3               (port1_P3),                                               //     .export
		.coe_P4               (port1_P4),                                               //     .export
		.coe_P5               (port1_P5),                                               //     .export
		.coe_P6               (port1_P6),                                               //     .export
		.coe_P7               (port1_P7)                                                //     .export
	);

	fan_motor_driver fan_motor_driver_0 (
		.rsi_MRST_reset       (qsys_serial_host_0_mrst_reset),                                      //      MRST.reset
		.csi_MCLK_clk         (qsys_serial_host_0_mclk_clk),                                        //      MCLK.clk
		.avs_ctrl_writedata   (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_writedata),   //      ctrl.writedata
		.avs_ctrl_readdata    (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_readdata),    //          .readdata
		.avs_ctrl_byteenable  (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_byteenable),  //          .byteenable
		.avs_ctrl_address     (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_address),     //          .address
		.avs_ctrl_write       (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_write),       //          .write
		.avs_ctrl_read        (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_read),        //          .read
		.avs_ctrl_waitrequest (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_waitrequest), //          .waitrequest
		.rsi_PWMRST_reset     (qsys_serial_host_0_mrst_reset),                                      //    PWMRST.reset
		.csi_PWMCLK_clk       (qsys_serial_host_0_mclk_clk),                                        //    PWMCLK.clk
		.fan                  (led_export)                                                          // fan_motor.export
	);

	fan_motor_driver fan_motor_driver_1 (
		.rsi_MRST_reset       (qsys_serial_host_0_mrst_reset),                                      //      MRST.reset
		.csi_MCLK_clk         (qsys_serial_host_0_mclk_clk),                                        //      MCLK.clk
		.avs_ctrl_writedata   (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_writedata),   //      ctrl.writedata
		.avs_ctrl_readdata    (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_readdata),    //          .readdata
		.avs_ctrl_byteenable  (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_byteenable),  //          .byteenable
		.avs_ctrl_address     (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_address),     //          .address
		.avs_ctrl_write       (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_write),       //          .write
		.avs_ctrl_read        (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_read),        //          .read
		.avs_ctrl_waitrequest (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_waitrequest), //          .waitrequest
		.rsi_PWMRST_reset     (qsys_serial_host_0_mrst_reset),                                      //    PWMRST.reset
		.csi_PWMCLK_clk       (qsys_serial_host_0_mclk_clk),                                        //    PWMCLK.clk
		.fan                  (humidifier_export)                                                   // fan_motor.export
	);

	fan_motor_driver fan_motor_driver_2 (
		.rsi_MRST_reset       (qsys_serial_host_0_mrst_reset),                                      //      MRST.reset
		.csi_MCLK_clk         (qsys_serial_host_0_mclk_clk),                                        //      MCLK.clk
		.avs_ctrl_writedata   (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_writedata),   //      ctrl.writedata
		.avs_ctrl_readdata    (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_readdata),    //          .readdata
		.avs_ctrl_byteenable  (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_byteenable),  //          .byteenable
		.avs_ctrl_address     (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_address),     //          .address
		.avs_ctrl_write       (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_write),       //          .write
		.avs_ctrl_read        (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_read),        //          .read
		.avs_ctrl_waitrequest (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_waitrequest), //          .waitrequest
		.rsi_PWMRST_reset     (qsys_serial_host_0_mrst_reset),                                      //    PWMRST.reset
		.csi_PWMCLK_clk       (qsys_serial_host_0_mclk_clk),                                        //    PWMCLK.clk
		.fan                  (humidifier_fan_export)                                               // fan_motor.export
	);

	brush_motor_driver brush_motor_driver_0 (
		.rsi_MRST_reset       (qsys_serial_host_0_mrst_reset),                                        //        MRST.reset
		.csi_MCLK_clk         (qsys_serial_host_0_mclk_clk),                                          //        MCLK.clk
		.avs_ctrl_writedata   (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_writedata),   //        ctrl.writedata
		.avs_ctrl_readdata    (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_readdata),    //            .readdata
		.avs_ctrl_byteenable  (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_byteenable),  //            .byteenable
		.avs_ctrl_address     (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_address),     //            .address
		.avs_ctrl_write       (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_write),       //            .write
		.avs_ctrl_read        (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_read),        //            .read
		.avs_ctrl_waitrequest (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_waitrequest), //            .waitrequest
		.HX                   (semi_cooler_HX),                                                       // brush_motor.export
		.HY                   (semi_cooler_HY),                                                       //            .export
		.rsi_PWMRST_reset     (qsys_serial_host_0_mrst_reset),                                        //      PWMRST.reset
		.csi_PWMCLK_clk       (qsys_serial_host_0_mclk_clk)                                           //      PWMCLK.clk
	);

	fan_motor_driver fan_motor_driver_3 (
		.rsi_MRST_reset       (qsys_serial_host_0_mrst_reset),                                      //      MRST.reset
		.csi_MCLK_clk         (qsys_serial_host_0_mclk_clk),                                        //      MCLK.clk
		.avs_ctrl_writedata   (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_writedata),   //      ctrl.writedata
		.avs_ctrl_readdata    (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_readdata),    //          .readdata
		.avs_ctrl_byteenable  (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_byteenable),  //          .byteenable
		.avs_ctrl_address     (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_address),     //          .address
		.avs_ctrl_write       (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_write),       //          .write
		.avs_ctrl_read        (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_read),        //          .read
		.avs_ctrl_waitrequest (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_waitrequest), //          .waitrequest
		.rsi_PWMRST_reset     (qsys_serial_host_0_mrst_reset),                                      //    PWMRST.reset
		.csi_PWMCLK_clk       (qsys_serial_host_0_mclk_clk),                                        //    PWMCLK.clk
		.fan                  (dryer_export)                                                        // fan_motor.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (8),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (0),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) qsys_serial_host_0_m1_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                              //                       clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                            //                     reset.reset
		.uav_address           (qsys_serial_host_0_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (qsys_serial_host_0_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (qsys_serial_host_0_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (qsys_serial_host_0_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (qsys_serial_host_0_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (qsys_serial_host_0_m1_byteenable),                                         //                          .byteenable
		.av_begintransfer      (qsys_serial_host_0_m1_begintransfer),                                      //                          .begintransfer
		.av_read               (qsys_serial_host_0_m1_read),                                               //                          .read
		.av_readdata           (qsys_serial_host_0_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (qsys_serial_host_0_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (qsys_serial_host_0_m1_write),                                              //                          .write
		.av_writedata          (qsys_serial_host_0_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                     //               (terminated)
		.av_chipselect         (1'b0),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                     //               (terminated)
		.av_debugaccess        (1'b0),                                                                     //               (terminated)
		.uav_clken             (),                                                                         //               (terminated)
		.av_clken              (1'b1)                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio8_0_gpio_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                            //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                          //                    reset.reset
		.uav_address           (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio8_0_gpio_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio8_0_gpio_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pio8_0_gpio_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pio8_0_gpio_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio8_0_gpio_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pio8_0_gpio_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (pio8_0_gpio_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio8_1_gpio_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                            //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                          //                    reset.reset
		.uav_address           (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio8_1_gpio_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio8_1_gpio_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pio8_1_gpio_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pio8_1_gpio_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio8_1_gpio_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pio8_1_gpio_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (pio8_1_gpio_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fan_motor_driver_0_ctrl_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                                        //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                                      //                    reset.reset
		.uav_address           (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (fan_motor_driver_0_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fan_motor_driver_1_ctrl_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                                        //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                                      //                    reset.reset
		.uav_address           (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (fan_motor_driver_1_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fan_motor_driver_2_ctrl_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                                        //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                                      //                    reset.reset
		.uav_address           (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (fan_motor_driver_2_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) brush_motor_driver_0_ctrl_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                                          //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                                        //                    reset.reset
		.uav_address           (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (brush_motor_driver_0_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_chipselect         (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fan_motor_driver_3_ctrl_translator (
		.clk                   (qsys_serial_host_0_mclk_clk),                                                        //                      clk.clk
		.reset                 (qsys_serial_host_0_mrst_reset),                                                      //                    reset.reset
		.uav_address           (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (fan_motor_driver_3_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_BEGIN_BURST           (65),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.PKT_BURST_TYPE_H          (62),
		.PKT_BURST_TYPE_L          (61),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_THREAD_ID_H           (73),
		.PKT_THREAD_ID_L           (73),
		.PKT_CACHE_H               (80),
		.PKT_CACHE_L               (77),
		.PKT_DATA_SIDEBAND_H       (64),
		.PKT_DATA_SIDEBAND_L       (64),
		.PKT_QOS_H                 (66),
		.PKT_QOS_L                 (66),
		.PKT_ADDR_SIDEBAND_H       (63),
		.PKT_ADDR_SIDEBAND_L       (63),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent (
		.clk              (qsys_serial_host_0_mclk_clk),                                                       //       clk.clk
		.reset            (qsys_serial_host_0_mrst_reset),                                                     // clk_reset.reset
		.av_address       (qsys_serial_host_0_m1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (qsys_serial_host_0_m1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (qsys_serial_host_0_m1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (qsys_serial_host_0_m1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (qsys_serial_host_0_m1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (qsys_serial_host_0_m1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (qsys_serial_host_0_m1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                             //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                              //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                              //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio8_0_gpio_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                      //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                    //       clk_reset.reset
		.m0_address              (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio8_0_gpio_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                      //                .channel
		.rf_sink_ready           (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                      //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                    // clk_reset.reset
		.in_data           (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio8_1_gpio_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                      //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                    //       clk_reset.reset
		.m0_address              (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio8_1_gpio_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                      //                .channel
		.rf_sink_ready           (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                      //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                    // clk_reset.reset
		.in_data           (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                                  //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                                //       clk_reset.reset
		.m0_address              (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                                  //                .channel
		.rf_sink_ready           (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                                  //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                                // clk_reset.reset
		.in_data           (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                                  //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                                //       clk_reset.reset
		.m0_address              (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                                  //                .channel
		.rf_sink_ready           (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                                  //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                                // clk_reset.reset
		.in_data           (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                                  //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                                //       clk_reset.reset
		.m0_address              (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src4_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_src4_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_src4_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_src4_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src4_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src4_channel),                                                                  //                .channel
		.rf_sink_ready           (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                                  //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                                // clk_reset.reset
		.in_data           (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                                    //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                                  //       clk_reset.reset
		.m0_address              (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src5_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_src5_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_src5_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_src5_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src5_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src5_channel),                                                                    //                .channel
		.rf_sink_ready           (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                                    //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                                  // clk_reset.reset
		.in_data           (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (65),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (57),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (60),
		.PKT_BURST_SIZE_L          (58),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (qsys_serial_host_0_mclk_clk),                                                                  //             clk.clk
		.reset                   (qsys_serial_host_0_mrst_reset),                                                                //       clk_reset.reset
		.m0_address              (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src6_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_src6_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_src6_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_src6_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src6_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src6_channel),                                                                  //                .channel
		.rf_sink_ready           (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (qsys_serial_host_0_mclk_clk),                                                                  //       clk.clk
		.reset             (qsys_serial_host_0_mrst_reset),                                                                // clk_reset.reset
		.in_data           (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	qsys_addr_router addr_router (
		.sink_ready         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (qsys_serial_host_0_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                       //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_src_valid),                                                             //          .valid
		.src_data           (addr_router_src_data),                                                              //          .data
		.src_channel        (addr_router_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                        //          .endofpacket
	);

	qsys_id_router id_router (
		.sink_ready         (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio8_0_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                            //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                          // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                    //       src.ready
		.src_valid          (id_router_src_valid),                                                    //          .valid
		.src_data           (id_router_src_data),                                                     //          .data
		.src_channel        (id_router_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                               //          .endofpacket
	);

	qsys_id_router id_router_001 (
		.sink_ready         (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio8_1_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                            //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                          // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                //       src.ready
		.src_valid          (id_router_001_src_valid),                                                //          .valid
		.src_data           (id_router_001_src_data),                                                 //          .data
		.src_channel        (id_router_001_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                           //          .endofpacket
	);

	qsys_id_router id_router_002 (
		.sink_ready         (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fan_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                        //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                            //       src.ready
		.src_valid          (id_router_002_src_valid),                                                            //          .valid
		.src_data           (id_router_002_src_data),                                                             //          .data
		.src_channel        (id_router_002_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                       //          .endofpacket
	);

	qsys_id_router id_router_003 (
		.sink_ready         (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fan_motor_driver_1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                        //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                            //       src.ready
		.src_valid          (id_router_003_src_valid),                                                            //          .valid
		.src_data           (id_router_003_src_data),                                                             //          .data
		.src_channel        (id_router_003_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                       //          .endofpacket
	);

	qsys_id_router id_router_004 (
		.sink_ready         (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fan_motor_driver_2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                        //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                            //       src.ready
		.src_valid          (id_router_004_src_valid),                                                            //          .valid
		.src_data           (id_router_004_src_data),                                                             //          .data
		.src_channel        (id_router_004_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                       //          .endofpacket
	);

	qsys_id_router id_router_005 (
		.sink_ready         (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (brush_motor_driver_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                          //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                              //       src.ready
		.src_valid          (id_router_005_src_valid),                                                              //          .valid
		.src_data           (id_router_005_src_data),                                                               //          .data
		.src_channel        (id_router_005_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                         //          .endofpacket
	);

	qsys_id_router id_router_006 (
		.sink_ready         (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fan_motor_driver_3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (qsys_serial_host_0_mclk_clk),                                                        //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                            //       src.ready
		.src_valid          (id_router_006_src_valid),                                                            //          .valid
		.src_data           (id_router_006_src_data),                                                             //          .data
		.src_channel        (id_router_006_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                       //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (70),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (7),
		.VALID_WIDTH               (7),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (qsys_serial_host_0_mclk_clk),    //       clk.clk
		.reset                  (qsys_serial_host_0_mrst_reset),  // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	qsys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (qsys_serial_host_0_mclk_clk),       //        clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),     //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_src6_endofpacket)    //           .endofpacket
	);

	qsys_rsp_xbar_demux rsp_xbar_demux (
		.clk                (qsys_serial_host_0_mclk_clk),       //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),     // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	qsys_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	qsys_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	qsys_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	qsys_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	qsys_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	qsys_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset              (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	qsys_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (qsys_serial_host_0_mclk_clk),           //       clk.clk
		.reset               (qsys_serial_host_0_mrst_reset),         // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

endmodule
